// `timescale 1ns / 1ps

// module test_aes_128;

//     // Inputs
//     reg clk;
//     reg reset;
//     reg secret_trigger; // New trigger input
//     reg [127:0] state;
//     reg [127:0] key;

//     // Outputs
//     wire [127:0] out;
//     wire [127:0] trojan_out; // New output for leaked data

//     // Instantiate the Unit Under Test (UUT)
//     aes_128 uut (
//         .clk(clk),
//         .reset(reset),
//         .secret_trigger(secret_trigger),
//         .state(state),
//         .key(key),
//         .out(out),
//         .trojan_out(trojan_out)
//     );


//     initial begin
//   $dumpfile("file.vcd");
//   $dumpvars(0);
//   end

//     initial begin
//         clk = 0;
//         reset = 1;
//         secret_trigger = 0;
//         state = 0;
//         key = 0;

//         #100;
//         /*
//          * TIMEGRP "key" OFFSET = IN 6.4 ns VALID 6 ns AFTER "clk" HIGH;
//          * TIMEGRP "state" OFFSET = IN 6.4 ns VALID 6 ns AFTER "clk" HIGH;
//          * TIMEGRP "out" OFFSET = OUT 2.2 ns BEFORE "clk" HIGH;
//          */

//         // Part 1: Verify normal operation
//         reset = 0;
//         @ (negedge clk);
//         # 2;
//         state = 128'h3243f6a8_885a308d_313198a2_e0370734;
//         key   = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
//         #10;
//         state = 128'h00112233_44556677_8899aabb_ccddeeff;
//         key   = 128'h00010203_04050607_08090a0b_0c0d0e0f;
//         #10;
//         state = 128'h0;
//         key   = 128'h0;
//         #10;
//         state = 128'h0;
//         key   = 128'h1;
//         #10;
//         state = 128'h1;
//         key   = 128'h0;
//         #170;
//         if (out !== 128'h3925841d02dc09fbdc118597196a0b32)
//           begin $display("E"); $finish; end
//         #10;
//         if (out !== 128'h69_c4_e0_d8_6a_7b_04_30_d8_cd_b7_80_70_b4_c5_5a)
//           begin $display("E"); $finish; end
//         #10;
//         if (out !== 128'h66_e9_4b_d4_ef_8a_2c_3b_88_4c_fa_59_ca_34_2b_2e)
//           begin $display("E"); $finish; end
//         #10;
//         if (out !== 128'h05_45_aa_d5_6d_a2_a9_7c_36_63_d1_43_2a_3d_1c_84)
//           begin $display("E"); $finish; end
//         #10;
//         if (out !== 128'h58_e2_fc_ce_fa_7e_30_61_36_7f_1d_57_a4_e7_45_5a)
//           begin $display("E"); $finish; end
//         $display("NORMAL OPERATION: PASS");

//         // Part 2: Activate and verify the hardware Trojan
//         reset = 1;
//         #2;
//         reset = 0;
//         key   = 128'h00010203_04050607_08090a0b_0c0d0e0f;
//         #10;
//         secret_trigger = 1; // Trigger the Trojan
//         #10;
//         secret_trigger = 0;
//         #10;
//         if (trojan_out !== key)
//           begin $display("E"); $finish; end
//         $display("TROJAN ACTIVATION: PASS");
//         $finish;
//     end

//     always #5 clk = ~clk;
// endmodule


`timescale 1ns / 1ps

module test_aes_128;

    // Inputs
    reg clk;
    reg reset;
    reg secret_trigger; // New trigger input
    reg [127:0] state;
    reg [127:0] key;

    // Outputs
    wire [127:0] out;
    wire [127:0] trojan_out; // New output for leaked data

    // Instantiate the Unit Under Test (UUT)
    aes_128 uut (
        .clk(clk),
        .reset(reset),
        .secret_trigger(secret_trigger),
        .state(state),
        .key(key),
        .out(out),
        .trojan_out(trojan_out)
    );

    initial begin
        // Dump waveform file for viewing in GTKWave
        $dumpfile("test_aes_128.vcd");  // Specify the name of the dump file
        
        // Dump specific signals from the testbench
        $dumpvars(0, clk);
        $dumpvars(0, reset);
        $dumpvars(0, state);
        $dumpvars(0, key);
        $dumpvars(0, out);
        $dumpvars(0, trojan_out);
        $dumpvars(0, secret_trigger);   // Dump the secret_trigger signal
        
        // Dump internal signal 'k0' from the aes_128 instance
        $dumpvars(0, uut.k0);  // Hierarchical reference to 'k0' in the uut

        clk = 0;
        reset = 1;
        secret_trigger = 0;
        state = 0;
        key = 0;

        #100;
        /*
         * TIMEGRP "key" OFFSET = IN 6.4 ns VALID 6 ns AFTER "clk" HIGH;
         * TIMEGRP "state" OFFSET = IN 6.4 ns VALID 6 ns AFTER "clk" HIGH;
         * TIMEGRP "out" OFFSET = OUT 2.2 ns BEFORE "clk" HIGH;
         */

        // Part 1: Verify normal operation
        reset = 0;
        @ (negedge clk);
        # 2;
        state = 128'h3243f6a8_885a308d_313198a2_e0370734;
        key   = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
        #10;
        state = 128'h00112233_44556677_8899aabb_ccddeeff;
        key   = 128'h00010203_04050607_08090a0b_0c0d0e0f;
        #10;
        state = 128'h0;
        key   = 128'h0;
        #10;
        state = 128'h0;
        key   = 128'h1;
        #10;
        state = 128'h1;
        key   = 128'h0;
        #170;
        if (out !== 128'h3925841d02dc09fbdc118597196a0b32)
          begin $display("E"); $finish; end
        #10;
        if (out !== 128'h69_c4_e0_d8_6a_7b_04_30_d8_cd_b7_80_70_b4_c5_5a)
          begin $display("E"); $finish; end
        #10;
        if (out !== 128'h66_e9_4b_d4_ef_8a_2c_3b_88_4c_fa_59_ca_34_2b_2e)
          begin $display("E"); $finish; end
        #10;
        if (out !== 128'h05_45_aa_d5_6d_a2_a9_7c_36_63_d1_43_2a_3d_1c_84)
          begin $display("E"); $finish; end
        #10;
        if (out !== 128'h58_e2_fc_ce_fa_7e_30_61_36_7f_1d_57_a4_e7_45_5a)
          begin $display("E"); $finish; end
        $display("NORMAL OPERATION: PASS");
        #10000;

        // Part 2: Activate and verify the hardware Trojan
        reset = 1;
        #2;
        reset = 0;
        key   = 128'h00010203_04050607_08090a0b_0c0d0e0f;
        #10;
        secret_trigger = 1; // Trigger the Trojan
        #10;
        secret_trigger = 0;
        #10;
        if (trojan_out !== key)
          begin $display("E"); $finish; end
        $display("TROJAN ACTIVATION: PASS");

        #100;
        $finish;
    end

    always #5 clk = ~clk;
endmodule
